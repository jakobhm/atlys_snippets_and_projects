--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package MAC_1G_RX_TYPES is

constant output_buffer_addr_width : integer := 4;
constant output_buffer_word_width : integer := 8;
constant output_buffer_addr_cnt   : integer := 15;

end MAC_1G_RX_TYPES;

package body MAC_1G_RX_TYPES is
 
end MAC_1G_RX_TYPES;
